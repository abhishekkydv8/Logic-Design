module and_gate(c,a,b);

output c;
input a,b;

wire x;

nand(x,a,b);
nand(c,x,x);

endmodule