module not_gate(b,a);

input a;
output b;

nand(b,a,a);

endmodule

