module not_gate(c,a,a);

output c;
input a;

nand(c,a,a);
endmodule
