module sub_16(diff,bout,in0,in1,bin);

output [15:0]diff;
output bout;

input [15:0]in0,in1;
input bin;

full_subtractor f1(diff[0],b0,in0[0],in1[0],bin);
full_subtractor f2(diff[1],b1,in0[1],in1[1],b0);
full_subtractor f3(diff[2],b2,in0[2],in1[2],b1);
full_subtractor f4(diff[3],b3,in0[3],in1[3],b2);

full_subtractor f5(diff[4],b4,in0[4],in1[4],b3);
full_subtractor f6(diff[5],b5,in0[5],in1[5],b4);
full_subtractor f7(diff[6],b6,in0[6],in1[6],b5);
full_subtractor f8(diff[7],b7,in0[7],in1[7],b6);

full_subtractor f9(diff[8],b8,in0[8],in1[8],b7);
full_subtractor f10(diff[9],b9,in0[9],in1[9],b8);
full_subtractor f11(diff[10],b10,in0[10],in1[10],b9);
full_subtractor f12(diff[11],b11,in0[11],in1[11],b10);

full_subtractor f13(diff[12],b12,in0[12],in1[12],b11);
full_subtractor f14(diff[13],b13,in0[13],in1[13],b12);
full_subtractor f15(diff[14],b14,in0[14],in1[14],b13);
full_subtractor f16(diff[15],bout,in0[15],in1[15],b14);

endmodule
