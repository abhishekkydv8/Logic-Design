module not_gate(a,b);
input b;
output a;
nand(a,b,b);
endmodule
 
