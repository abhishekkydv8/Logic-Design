module not16_gate(b,a);

output[15:0]b;
input[15:0]a;

not_gate not_gate_16[15:0](b,a);

endmodule

